LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
ENTITY NiosFighter IS
PORT (
		SW : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		KEY : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CLOCK_50 : IN STD_LOGIC;
		LEDG : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		DRAM_CLK, DRAM_CKE : OUT STD_LOGIC;
		DRAM_ADDR : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
		DRAM_BA_0, DRAM_BA_1 : BUFFER STD_LOGIC;
		DRAM_CS_N, DRAM_CAS_N, DRAM_RAS_N, DRAM_WE_N : OUT STD_LOGIC;
		DRAM_DQ : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		DRAM_UDQM, DRAM_LDQM : BUFFER STD_LOGIC;
		LCD_DATA : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		LCD_ON, LCD_BLON, LCD_EN, LCD_RS, LCD_RW : OUT STD_LOGIC;
		VGA_R, VGA_G, VGA_B : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		VGA_CLK, VGA_BLANK, VGA_HS,VGA_VS, VGA_SYNC : OUT STD_LOGIC;
		SRAM_DQ: INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		SRAM_ADDR: OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
		SRAM_LB_N, SRAM_UB_N,SRAM_CE_N,SRAM_OE_N,SRAM_WE_N: OUT STD_LOGIC;
		SD_CMD : inout std_logic;
		SD_DAT : inout std_logic;
		SD_DAT3: inout std_logic;
		SD_CLK : out   std_logic;
		I2C_SCLK: out   std_logic;
		I2C_SDAT:inout std_logic);
END NiosFighter;
ARCHITECTURE Structure OF NiosFighter IS
COMPONENT fighterSystem
PORT (
		clk_clk : IN STD_LOGIC;
		reset_reset_n : IN STD_LOGIC;
		sdram_clk_clk : OUT STD_LOGIC;
		leds_export : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		switches_export : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		sdram_wire_addr : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
		sdram_wire_ba : BUFFER STD_LOGIC_VECTOR(1 DOWNTO 0);
		sdram_wire_cas_n : OUT STD_LOGIC;
		sdram_wire_cke : OUT STD_LOGIC;
		sdram_wire_cs_n : OUT STD_LOGIC;
		sdram_wire_dq : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		sdram_wire_dqm : BUFFER STD_LOGIC_VECTOR(1 DOWNTO 0);
		sdram_wire_ras_n : OUT STD_LOGIC;
		sdram_wire_we_n : OUT STD_LOGIC;
		lcd_data_DATA : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		lcd_data_ON : OUT STD_LOGIC;
		lcd_data_BLON : OUT STD_LOGIC;
		lcd_data_EN : OUT STD_LOGIC;
		lcd_data_RS : OUT STD_LOGIC;
		lcd_data_RW : OUT STD_LOGIC;
		vga_controller_R : OUT std_logic_vector(9 DOWNTO 0);
		vga_controller_G : OUT std_logic_vector(9 DOWNTO 0);
		vga_controller_B : OUT std_logic_vector(9 DOWNTO 0);
		vga_controller_CLK : OUT std_logic;
		vga_controller_BLANK : OUT std_logic;
		vga_controller_HS : OUT std_logic;
		vga_controller_VS : OUT std_logic;
		vga_controller_SYNC:OUT std_logic;
		SRAM_DQ : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		SRAM_ADDR : OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
		SRAM_LB_N : OUT STD_LOGIC;
		SRAM_UB_N : OUT STD_LOGIC;
		SRAM_CE_N : OUT STD_LOGIC;
		SRAM_OE_N : OUT STD_LOGIC;
		SRAM_WE_N : OUT STD_LOGIC;
		key_export : in std_logic_vector(3 downto 0);
		sd_card_b_SD_cmd     : inout std_logic;
		sd_card_b_SD_dat     : inout std_logic;
		sd_card_b_SD_dat3    : inout std_logic;
		sd_card_o_SD_clock   : out   std_logic;
		audio_SDAT           : inout std_logic;
      audio_SCLK           : out   std_logic );
END COMPONENT;
SIGNAL DQM : STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL BA : STD_LOGIC_VECTOR(1 DOWNTO 0);
BEGIN
DRAM_BA_0<= BA(0);
DRAM_BA_1<= BA(1);
DRAM_UDQM<= DQM(1);
DRAM_LDQM<= DQM(0);
--Instantiate the Nios II system entity generated by the Qsys tool.
NiosII: fighterSystem
PORT MAP (
		clk_clk => CLOCK_50,
		reset_reset_n => SW(1),
		sdram_clk_clk => DRAM_CLK,
		leds_export => LEDG,
		switches_export => SW,
		sdram_wire_addr => DRAM_ADDR,
		sdram_wire_ba => BA,
		sdram_wire_cas_n => DRAM_CAS_N,
		sdram_wire_cke => DRAM_CKE,
		sdram_wire_cs_n => DRAM_CS_N,
		sdram_wire_dq => DRAM_DQ,
		sdram_wire_dqm => DQM,
		sdram_wire_ras_n => DRAM_RAS_N,
		sdram_wire_we_n => DRAM_WE_N,
		lcd_data_DATA => LCD_DATA,
		lcd_data_ON => LCD_ON,
		lcd_data_BLON => LCD_BLON,
		lcd_data_EN => LCD_EN,
		lcd_data_RS => LCD_RS,
		lcd_data_RW => LCD_RW,
		vga_controller_CLK => VGA_CLK,
		vga_controller_HS => VGA_HS,
		vga_controller_VS => VGA_VS,
		vga_controller_BLANK => VGA_BLANK,
		vga_controller_SYNC => VGA_SYNC,
		vga_controller_R => VGA_R,
		vga_controller_G => VGA_G,
		vga_controller_B => VGA_B,
		sram_DQ => SRAM_DQ,
		sram_ADDR => SRAM_ADDR,
		sram_LB_N => SRAM_LB_N,
		sram_UB_N => SRAM_UB_N,
		sram_CE_N => SRAM_CE_N,
		sram_OE_N => SRAM_OE_N,
		sram_WE_N => SRAM_WE_N,
		key_export => KEY,
		sd_card_b_SD_cmd     => SD_CMD,
		sd_card_b_SD_dat     => SD_DAT,
		sd_card_b_SD_dat3    => SD_DAT3,
		sd_card_o_SD_clock   => SD_CLK,
		audio_SDAT =>I2C_SDAT,
      audio_SCLK =>I2C_SCLK);
END Structure;