--NiosFighter.vhdl