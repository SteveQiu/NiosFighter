--TEst2